`timescale 1ps/1ps

module simonEncyrpt_tb;
		parameter WIDTH = 64;
		parameter size = 46875; //#rows of file - look it up because Verilog doesnt recognize $size()
		reg [63:0] A [0:size-1];
		integer f_out,i;
		reg [63:0] indata  = 64'b1011101000111010001110100011101000111011001110110011110000111100;
		wire [127:0] keySeedval = 128'b10110100011111101000111001011001011111100010110101010100111101000100100110101100100001010101111101010101011000101111010011100111;
		//10110100011111101000111001011001011111100010110101010100111101000100100110101100100001010101111101010101011000101111010011100111
		//11111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111111
		//00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000
		//00000000000000000000000000000000000000000000000000000000000000001111111111111111111111111111111111111111111111111111111111111111
		wire [63:0] outvalue;
		simonEncrypt encrypt1 (.input_Val(indata), .keySeed(keySeedval), .encrypted_Val(outvalue));

	initial begin
		$readmemb("complex_64b_binary.txt",A);
		//f_out = $fopen("bin_encrypt_complex.txt","w");
		//f_out = $fopen("roundKeys_simple2.txt","w");

		for (i = 0; i<size; i=i+1) begin
			//indata = A[i];
			#1;
			$display("i=%d: indata=%b outdata=%b #remaining:%d",i,indata,outvalue,size-1-i);
			//$fdisplay(f_out,"%b",outvalue);
		end
		//$fclose(f_out);
		//$stop;
	end
endmodule

